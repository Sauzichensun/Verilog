module moduleName (
    input wire clk,
    input wire rst,
    output wire [7:0] data_out
);
endmodule

