module teset (
    input a,
    output b
);
    assign b = a;
endmodule

